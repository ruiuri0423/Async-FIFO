// Including all sub-module
//--------------------------------
`include "CNT_empty.v"
`include "CNT_full.v"
`include "DFF.v"
`include "DFF_n.v"
`include "RF.v"
`include "Synchronizer.v"
//--------------------------------
// End